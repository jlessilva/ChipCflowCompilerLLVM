decider x,y,zforicexx x1,x2,x3,x4,x5; 
add x1,x2,x3; 
